module area(
   input [8:0] ax,
   input [8:0] bx,
   input [8:0] cx,
   input [8:0] ay,
   input [8:0] by,
   input [8:0] cy,
   output [17:0] area
);

always @( ax or bx .. ) 

// 

endmodule
