module testbench;



endmodule
